library IEEE;
use IEEE.Std_logic_1164.all;
use IEEE.Numeric_Std.all;

entity SigmaDeltaConverter is
  
end entity SigmaDeltaConverter;

architecture code of SigmaDeltaConverter is
  
begin
  
  
  
  
  
end architecture;
